
----------------------------------------------------------------
-- Instruction Memory
----------------------------------------------------------------
constant INSTR_MEM : MEM_128x32 := (		x"EB000040", 
											x"E480D000", 
											x"EB000041", 
											x"E480D001", 
											x"E3A03001", 
											x"E3A09003", 
											x"E3A0A801", 
											x"E24AA001", 
											x"E59F81D8", 
											x"E1A00000", 
											x"E5980004", 
											x"E0101913", 
											x"0AFFFFFC", 
											x"E5984000", 
											x"E004400A", 
											x"E5980004", 
											x"E0101183", 
											x"1AFFFFFC", 
											x"E5980004", 
											x"E0101913", 
											x"0AFFFFFC", 
											x"E5985000", 
											x"E2055007", 
											x"E5980004", 
											x"E0101183", 
											x"1AFFFFFC", 
											x"E5980004", 
											x"E0101913", 
											x"0AFFFFFC", 
											x"E5986000", 
											x"E006600A", 
											x"E5980004", 
											x"E0101183", 
											x"1AFFFFFC", 
											x"E3550000", 
											x"0A00000C", 
											x"E3550001", 
											x"0A00000C", 
											x"E3550002", 
											x"0A00000C", 
											x"E3550003", 
											x"0A00000C", 
											x"E3350004", 
											x"0A00000C", 
											x"E3350005", 
											x"0A00000C", 
											x"E3350006", 
											x"0A00000C", 
											x"1A00000D", 
											x"E0847006", 
											x"EA00000C", 
											x"E0447006", 
											x"EA00000A", 
											x"E0070694", 
											x"EA000008", 
											x"E0275694", 
											x"EA000006", 
											x"E1C47006", 
											x"EA000004", 
											x"E0247006", 
											x"EA000002", 
											x"E0647006", 
											x"EA000000", 
											x"E0C47006", 
											x"E5087004", 
											x"EAFFFFC7", 
											x"E59FB0F4", 
											x"E588B014", 
											x"E1A0F00E", 
											x"E59FB0EC", 
											x"E588B014", 
											x"E1A0F00E", 
											others => x"00000000");

----------------------------------------------------------------
-- Data (Constant) Memory
----------------------------------------------------------------
constant DATA_CONST_MEM : MEM_128x32 := (	x"00000C04", 
											x"00002215", 
											x"22150000", 
											others => x"00000000");

